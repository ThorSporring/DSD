library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity my_and is
	
	port
	(
		-- Input ports
		a,b: in  std_logic;
		
		-- Output ports
		f	: out std_logic
	);
end my_and;

architecture my_and_impl of my_and is

begin
	f <= a and b;
end my_and_impl;


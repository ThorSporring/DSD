library verilog;
use verilog.vl_types.all;
entity meemoo_tester_vlg_vec_tst is
end meemoo_tester_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity code_lock_simple_vlg_vec_tst is
end code_lock_simple_vlg_vec_tst;
